library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity tubes2 is
port (y:out std_logic_vector(0 downto 255));

end entity;

architecture arch_tubes2 of tubes2 is
begin
	y<="0000000000000000000000000000000011111111000000000000000000000000000000001111111100000000000000000000010000000100111111110000010000000100000001000000010011111111000001000000010000000100000001001111111100011100001111000011110000011000";
		

end architecture; 